// CDLFont.cdl

Name: CDL Font
Version: 1.0
UID: 0x102045DC
Flag: KCdlFlagRomOnly

%% C++

#include <CdlFont.h>

%% API

TCdlArray<SIdMetricsPair> metricsArray;
TCdlArray<SLogicalIdMetricsIdPair> logicalIdMapArray;
