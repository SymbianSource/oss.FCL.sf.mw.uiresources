// This CDL file contains all excluded layout APIs

Name: Excluded
Version: 1.0
UID: 0x00000000

%% API

TAknLayoutTableLimits Grid_pane_descendants_SUB_TABLE_1_Limits();
TAknWindowLineLayout Grid_pane_descendants_SUB_TABLE_1(TInt aLineIndex, TInt aIndex_l, TInt aIndex_t);
TAknLayoutTableLimits Presence_status_list_components_Limits();
TAknWindowLineLayout Presence_status_list_components(TInt aLineIndex);
TAknLayoutTableLimits IM_chat_view_descendant_panes_Limits();
TAknWindowLineLayout IM_chat_view_descendant_panes(TInt aLineIndex, TInt aCommon1);
TAknLayoutTableLimits Media_Player_Playback_view_elements_Limits();
TAknWindowLineLayout Media_Player_Playback_view_elements(TInt aLineIndex);
TAknLayoutTableLimits SMIL_text_pane_elements_Limits();
TAknWindowLineLayout SMIL_text_pane_elements(TInt aLineIndex, const TRect& aParentRect);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_0_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_1_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_1(TInt aLineIndex);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_2_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_2(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_3_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_3(TInt aLineIndex);
TAknLayoutTableLimits Additional_heading_pane_elements_Limits();
TAknWindowLineLayout Additional_heading_pane_elements(TInt aLineIndex);
TAknWindowLineLayout scroll_pane(TInt aIndex_H); // excluded disallowed generated API name (duplicate lines same name) but only appears once in a variant
TAknLayoutTableLimits Message_writing_layout_elements_SUB_TABLE_0_Limits();
TAknWindowLineLayout Message_writing_layout_elements_SUB_TABLE_0(TInt aLineIndex, TInt aIndex_t, TInt aIndex_H);
TAknLayoutTableLimits Calendar_Week_view_elements_SUB_TABLE_1_Limits();
TAknWindowLineLayout Calendar_Week_view_elements_SUB_TABLE_1(TInt aLineIndex, TInt aIndex_t);
TAknLayoutTableLimits Pinboard_elements__list__SUB_TABLE_1_Limits();
TAknWindowLineLayout Pinboard_elements__list__SUB_TABLE_1(TInt aLineIndex);
TAknLayoutTableLimits IM_chat_view_descendant_panes_SUB_TABLE_0_Limits();
TAknWindowLineLayout IM_chat_view_descendant_panes_SUB_TABLE_0(TInt aLineIndex, TInt aCommon1);
TAknWindowLineLayout Presence_status_popup_window_elements_Line_1();
TAknLayoutTableLimits Calendar_Week_view_elements_SUB_TABLE_2_Limits();
TAknWindowLineLayout Calendar_Week_view_elements_SUB_TABLE_2(TInt aLineIndex);
