// This CDL file contains all excluded layout APIs

Name: Excluded
Version: 1.0
UID: 0x00000000

%% API

TAknLayoutTableLimits Status_pane_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Status_pane_descendants_SUB_TABLE_0(TInt aLineIndex, const TRect& aParentRect);
TAknLayoutTableLimits Navi_pane_texts_SUB_TABLE_0_Limits();
TAknTextLineLayout Navi_pane_texts_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Main_pane_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Main_pane_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknWindowLineLayout List_pane_elements__double_large_graphic__Line_11(TInt aIndex_l);
TAknLayoutTableLimits Form_pop_up_field_elements_and_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_pop_up_field_elements_and_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Form_pop_up_wide_field_elements_and_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_pop_up_wide_field_elements_and_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Form_slider_field_elements_and_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_slider_field_elements_and_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Form_slider_field_elements_and_descendants_dup_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_slider_field_elements_and_descendants_dup_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits List_pane_elements_and_descendants__settings_edited__SUB_TABLE_0_Limits();
TAknWindowLineLayout List_pane_elements_and_descendants__settings_edited__SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits List_pane_elements_and_descendants__settings_edited__SUB_TABLE_1_Limits();
TAknWindowLineLayout List_pane_elements_and_descendants__settings_edited__SUB_TABLE_1(TInt aLineIndex);
TAknLayoutTableLimits Pop_up_window_list_pane_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Pop_up_window_list_pane_descendants_SUB_TABLE_0(TInt aLineIndex, TInt aIndex_t);
TAknLayoutTableLimits List_pane_elements__menu_single_graphic_heading__SUB_TABLE_0_Limits();
TAknWindowLineLayout List_pane_elements__menu_single_graphic_heading__SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Data_query_pop_up_window_elements_SUB_TABLE_0_Limits();
TAknWindowLineLayout Data_query_pop_up_window_elements_SUB_TABLE_0(TInt aLineIndex, const TRect& aParentRect, TInt aCommon1);
TAknLayoutTableLimits Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_0_Limits();
TAknWindowLineLayout Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_0(TInt aLineIndex, TInt aIndex_C, TInt aIndex_t);
TAknLayoutTableLimits Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_1_Limits();
TAknWindowLineLayout Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_1(TInt aLineIndex, TInt aIndex_t);
TAknLayoutTableLimits Colour_selection_pop_up_window_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Colour_selection_pop_up_window_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits List_pane_elements__double_large_graphic__SUB_TABLE_0_Limits();
TAknWindowLineLayout List_pane_elements__double_large_graphic__SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_0_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_0(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_1_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_1(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_2_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_2(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Main_pane_descendants_SUB_TABLE_1_Limits();
TAknWindowLineLayout Main_pane_descendants_SUB_TABLE_1(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Grid_pane_descendants_SUB_TABLE_1_Limits();
TAknWindowLineLayout Grid_pane_descendants_SUB_TABLE_1(TInt aLineIndex, TInt aIndex_l, TInt aIndex_t);
TAknLayoutTableLimits Presence_status_list_components_Limits();
TAknWindowLineLayout Presence_status_list_components(TInt aLineIndex);
TAknLayoutTableLimits IM_chat_view_descendant_panes_Limits();
TAknWindowLineLayout IM_chat_view_descendant_panes(TInt aLineIndex, TInt aCommon1);
TAknLayoutTableLimits Media_Player_Playback_view_elements_Limits();
TAknWindowLineLayout Media_Player_Playback_view_elements(TInt aLineIndex);
TAknLayoutTableLimits SMIL_text_pane_elements_Limits();
TAknWindowLineLayout SMIL_text_pane_elements(TInt aLineIndex, const TRect& aParentRect);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_3_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_3(TInt aLineIndex);
TAknLayoutTableLimits Additional_heading_pane_elements_Limits();
TAknWindowLineLayout Additional_heading_pane_elements(TInt aLineIndex);

