// This CDL file contains all excluded layout APIs

Name: Excluded
Version: 1.0
UID: 0x00000000

%% API

TAknLayoutTableLimits Status_pane_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Status_pane_descendants_SUB_TABLE_0(TInt aLineIndex, const TRect& aParentRect);
TAknLayoutTableLimits Navi_pane_texts_SUB_TABLE_0_Limits();
TAknTextLineLayout Navi_pane_texts_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Main_pane_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Main_pane_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknWindowLineLayout List_pane_elements__double_large_graphic__Line_11(TInt aIndex_l);
TAknLayoutTableLimits Form_pop_up_field_elements_and_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_pop_up_field_elements_and_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknWindowLineLayout Form_pop_up_field_elements_and_descendants_SUB_TABLE_0(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Form_pop_up_wide_field_elements_and_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_pop_up_wide_field_elements_and_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Form_slider_field_elements_and_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_slider_field_elements_and_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Form_slider_field_elements_and_descendants_dup_SUB_TABLE_0_Limits();
TAknWindowLineLayout Form_slider_field_elements_and_descendants_dup_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits List_pane_elements_and_descendants__settings_edited__SUB_TABLE_0_Limits();
TAknWindowLineLayout List_pane_elements_and_descendants__settings_edited__SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits List_pane_elements_and_descendants__settings_edited__SUB_TABLE_1_Limits();
TAknWindowLineLayout List_pane_elements_and_descendants__settings_edited__SUB_TABLE_1(TInt aLineIndex);
TAknLayoutTableLimits Pop_up_window_list_pane_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Pop_up_window_list_pane_descendants_SUB_TABLE_0(TInt aLineIndex, TInt aIndex_t);
TAknLayoutTableLimits List_pane_elements__menu_single_graphic_heading__SUB_TABLE_0_Limits();
TAknWindowLineLayout List_pane_elements__menu_single_graphic_heading__SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Data_query_pop_up_window_elements_SUB_TABLE_0_Limits();
TAknWindowLineLayout Data_query_pop_up_window_elements_SUB_TABLE_0(TInt aLineIndex, const TRect& aParentRect, TInt aCommon1);
TAknLayoutTableLimits Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_0_Limits();
TAknWindowLineLayout Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_0(TInt aLineIndex, TInt aIndex_C, TInt aIndex_t);
TAknLayoutTableLimits Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_1_Limits();
TAknWindowLineLayout Combined_data_and_code_query_pop_up_window_elements_SUB_TABLE_1(TInt aLineIndex, TInt aIndex_t);
TAknLayoutTableLimits Colour_selection_pop_up_window_descendants_SUB_TABLE_0_Limits();
TAknWindowLineLayout Colour_selection_pop_up_window_descendants_SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits List_pane_elements__double_large_graphic__SUB_TABLE_0_Limits();
TAknWindowLineLayout List_pane_elements__double_large_graphic__SUB_TABLE_0(TInt aLineIndex);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_0_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_0(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_1_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_1(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_2_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_2(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Main_pane_descendants_SUB_TABLE_1_Limits();
TAknWindowLineLayout Main_pane_descendants_SUB_TABLE_1(TInt aLineIndex, TInt aIndex_H);
TAknLayoutTableLimits Pop_up_windows__main_pane_as_parent__SUB_TABLE_3_Limits();
TAknWindowLineLayout Pop_up_windows__main_pane_as_parent__SUB_TABLE_3(TInt aLineIndex);
TAknWindowLineLayout slider_set_pane(); // excluded disallowed generated API name (duplicate lines same name) but only appears once in a variant
TAknWindowLineLayout popup_submenu_window(TInt aCommon1); // excluded disallowed generated API name (duplicate lines same name) but only appears once in a variant
TAknWindowLineLayout scroll_pane(TInt aIndex_H); // excluded disallowed generated API name (duplicate lines same name) but only appears once in a variant
TAknLayoutTableLimits Fast_application_swapping_pop_up_window_graphics_Limits();
TAknWindowLineLayout Fast_application_swapping_pop_up_window_graphics(TInt aLineIndex, const TRect& aParentRect);
